module high_bit_search(
    input clk,
    input signed [INPUT_WIDTH-1:0] input_data,

    output reg signed [RESULT_WIDTH-1:0]result = 0
);

endmodule